LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY DivisorDeFrecuencia IS
	PORT (
		CLK100MHZ : IN STD_LOGIC;
		CLK : OUT STD_LOGIC
	);

END DivisorDeFrecuencia;
ARCHITECTURE Arquitectura OF DivisorDeFrecuencia IS
	CONSTANT MAX_COUNT : INTEGER := 50000000;
	SIGNAL COUNT : INTEGER RANGE 0 TO MAX_COUNT;
	SIGNAL CLK_STATE : STD_LOGIC := '0';

BEGIN
	GEN_CLOCK : PROCESS (CLK100MHZ, CLK_STATE, COUNT)
	BEGIN
		IF CLK100MHZ'EVENT AND CLK100MHZ = '1' THEN
			IF COUNT < MAX_COUNT THEN
 				COUNT <= COUNT + 1;
 			ELSE
 				CLK_STATE <= NOT CLK_STATE;
 				COUNT <= 0;
 			END IF;
 		END IF;
	END PROCESS;
	PERSECOND : PROCESS (CLK_STATE)
	BEGIN
		CLK <= CLK_STATE;
 	END PROCESS;
 END Arquitectura;